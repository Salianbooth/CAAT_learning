LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY RF IS
 PORT (
 CO :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 C0 :OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
 C1 : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
 C2 : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
 C3 : OUT STD_LOGIC_VECTOR(0 DOWNTO 0) );
END RF;
ARCHITECTURE behav OF RF IS
--SIGNAL OP : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
-- OP <= OP3&OP2&OP1&OP0;
 PROCESS(CO)
 BEGIN
 CASE CO IS
 WHEN "00"=> C0<="1";C1<="0";C2<="0";C3<="0";
 WHEN "01"=> C0<="0";C1<="1";C2<="0";C3<="0";
 WHEN "10"=> C0<="0";C1<="0";C2<="1";C3<="0";
 WHEN "11"=> C0<="0";C1<="0";C2<="0";C3<="1";
 END CASE;
 END PROCESS;
END behav;