-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Full Version"
-- CREATED		"Mon Jun 05 15:42:46 2023"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY computer IS 
	PORT
	(
		clock :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		ALUOUT1 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		ALUOUT2 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		ALUOUT3 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		ALUOUT4 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		s :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END computer;

ARCHITECTURE bdf_type OF computer IS 

COMPONENT alu_8b
	PORT(A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 S : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CO : OUT STD_LOGIC;
		 ZF : OUT STD_LOGIC;
		 F : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ram0
	PORT(wren : IN STD_LOGIC;
		 rden : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT data_mux
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT rf
	PORT(CO : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 C0 : OUT STD_LOGIC_VECTOR(0 TO 0);
		 C1 : OUT STD_LOGIC_VECTOR(0 TO 0);
		 C2 : OUT STD_LOGIC_VECTOR(0 TO 0);
		 C3 : OUT STD_LOGIC_VECTOR(0 TO 0)
	);
END COMPONENT;

COMPONENT ac_a
	PORT(LOAD_A : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 Data_in : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 A : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT immediate_mux
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux1
	PORT(data0x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT seg7_16b
	PORT(Blank : IN STD_LOGIC;
		 Test : IN STD_LOGIC;
		 Data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 RQ1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 RQ2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT rinstructiondecoder
	PORT(OP : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_constant0
	PORT(		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT controlunit
	PORT(OP : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 beq : OUT STD_LOGIC_VECTOR(0 TO 0);
		 bgt : OUT STD_LOGIC_VECTOR(0 TO 0);
		 bne : OUT STD_LOGIC_VECTOR(0 TO 0);
		 Exop : OUT STD_LOGIC_VECTOR(0 TO 0);
		 Imux1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 jump : OUT STD_LOGIC_VECTOR(0 TO 0);
		 ld : OUT STD_LOGIC_VECTOR(0 TO 0);
		 Lmux : OUT STD_LOGIC_VECTOR(0 TO 0);
		 PC_1 : OUT STD_LOGIC_VECTOR(0 TO 0);
		 R_tybe : OUT STD_LOGIC_VECTOR(0 TO 0);
		 S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Smux : OUT STD_LOGIC_VECTOR(0 TO 0);
		 str : OUT STD_LOGIC_VECTOR(0 TO 0);
		 WE : OUT STD_LOGIC_VECTOR(0 TO 0);
		 wpc : OUT STD_LOGIC_VECTOR(0 TO 0)
	);
END COMPONENT;

COMPONENT bit_mux
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pc
	PORT(clk : IN STD_LOGIC;
		 Reset : IN STD_LOGIC;
		 LOAD_PC : IN STD_LOGIC;
		 INCR_PC : IN STD_LOGIC;
		 Addr_Val_in : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 PC_out : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT offset
	PORT(in_c : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 out_c : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT address
	PORT(in_c : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 out_c : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_constant1
	PORT(		 result : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT immediate
	PORT(in_c : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 went : IN STD_LOGIC_VECTOR(0 TO 0);
		 out_c : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT adder_16bit
	PORT(A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 CarryOut : OUT STD_LOGIC;
		 Sum : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT rom0
	PORT(clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux0
	PORT(sel : IN STD_LOGIC;
		 data0x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	beq :  STD_LOGIC;
SIGNAL	bgt :  STD_LOGIC;
SIGNAL	bne :  STD_LOGIC;
SIGNAL	CO :  STD_LOGIC;
SIGNAL	DATA_A :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	DATA_B :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	exop :  STD_LOGIC;
SIGNAL	HALT :  STD_LOGIC;
SIGNAL	INCR_PC :  STD_LOGIC;
SIGNAL	IY_OUT :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	LMUX :  STD_LOGIC;
SIGNAL	LOAD_PC :  STD_LOGIC;
SIGNAL	PC_OUT :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	R_TY :  STD_LOGIC;
SIGNAL	WE :  STD_LOGIC;
SIGNAL	wpc :  STD_LOGIC;
SIGNAL	WRITE :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	WRITE_0 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	WRITE_1 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	ZF :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(3 DOWNTO 0);


BEGIN 
s <= SYNTHESIZED_WIRE_2;
SYNTHESIZED_WIRE_51 <= '0';
SYNTHESIZED_WIRE_52 <= '1';



SYNTHESIZED_WIRE_8 <= WE AND SYNTHESIZED_WIRE_0;


b2v_inst10 : alu_8b
PORT MAP(A => DATA_A,
		 B => SYNTHESIZED_WIRE_1,
		 S => SYNTHESIZED_WIRE_2,
		 CO => CO,
		 ZF => ZF,
		 F => WRITE_0);


b2v_inst12 : ram0
PORT MAP(wren => SYNTHESIZED_WIRE_3,
		 rden => WE,
		 clock => clock,
		 address => WRITE_0,
		 data => DATA_B,
		 q => WRITE_1);


SYNTHESIZED_WIRE_3 <= NOT(WE);



b2v_inst14 : data_mux
PORT MAP(sel => LMUX,
		 data0x => WRITE_0,
		 data1x => WRITE_1,
		 result => WRITE);


b2v_inst15 : rf
PORT MAP(CO => SYNTHESIZED_WIRE_4,
		 C0(0) => SYNTHESIZED_WIRE_0,
		 C1(0) => SYNTHESIZED_WIRE_5,
		 C2(0) => SYNTHESIZED_WIRE_6,
		 C3(0) => SYNTHESIZED_WIRE_7);


SYNTHESIZED_WIRE_10 <= WE AND SYNTHESIZED_WIRE_5;


SYNTHESIZED_WIRE_11 <= WE AND SYNTHESIZED_WIRE_6;


SYNTHESIZED_WIRE_12 <= WE AND SYNTHESIZED_WIRE_7;


b2v_inst19 : ac_a
PORT MAP(LOAD_A => SYNTHESIZED_WIRE_8,
		 clk => clock,
		 Data_in => WRITE,
		 A => SYNTHESIZED_WIRE_47);


b2v_inst2 : immediate_mux
PORT MAP(sel => R_TY,
		 data0x => DATA_B,
		 data1x => SYNTHESIZED_WIRE_9,
		 result => SYNTHESIZED_WIRE_1);


b2v_inst20 : ac_a
PORT MAP(LOAD_A => SYNTHESIZED_WIRE_10,
		 clk => clock,
		 Data_in => WRITE,
		 A => SYNTHESIZED_WIRE_48);


b2v_inst21 : ac_a
PORT MAP(LOAD_A => SYNTHESIZED_WIRE_11,
		 clk => clock,
		 Data_in => WRITE,
		 A => SYNTHESIZED_WIRE_49);


b2v_inst22 : ac_a
PORT MAP(LOAD_A => SYNTHESIZED_WIRE_12,
		 clk => clock,
		 Data_in => WRITE,
		 A => SYNTHESIZED_WIRE_50);


b2v_inst23 : lpm_mux1
PORT MAP(data0x => SYNTHESIZED_WIRE_47,
		 data1x => SYNTHESIZED_WIRE_48,
		 data2x => SYNTHESIZED_WIRE_49,
		 data3x => SYNTHESIZED_WIRE_50,
		 sel => IY_OUT(11 DOWNTO 10),
		 result => DATA_A);


b2v_inst24 : lpm_mux1
PORT MAP(data0x => SYNTHESIZED_WIRE_47,
		 data1x => SYNTHESIZED_WIRE_48,
		 data2x => SYNTHESIZED_WIRE_49,
		 data3x => SYNTHESIZED_WIRE_50,
		 sel => IY_OUT(9 DOWNTO 8),
		 result => DATA_B);


b2v_inst25 : seg7_16b
PORT MAP(Blank => SYNTHESIZED_WIRE_51,
		 Test => SYNTHESIZED_WIRE_52,
		 Data => WRITE_0(7 DOWNTO 0),
		 RQ1 => ALUOUT1,
		 RQ2 => ALUOUT2);


b2v_inst26 : seg7_16b
PORT MAP(Blank => SYNTHESIZED_WIRE_51,
		 Test => SYNTHESIZED_WIRE_52,
		 Data => WRITE_0(15 DOWNTO 8),
		 RQ1 => ALUOUT3,
		 RQ2 => ALUOUT4);



b2v_inst3 : rinstructiondecoder
PORT MAP(OP => IY_OUT(2 DOWNTO 0),
		 S => SYNTHESIZED_WIRE_45);


b2v_inst30 : data_mux
PORT MAP(sel => SYNTHESIZED_WIRE_25,
		 data0x => SYNTHESIZED_WIRE_53,
		 data1x => SYNTHESIZED_WIRE_27,
		 result => SYNTHESIZED_WIRE_28);


b2v_inst31 : lpm_constant0
PORT MAP(		 result => SYNTHESIZED_WIRE_43);


b2v_inst32 : data_mux
PORT MAP(sel => LOAD_PC,
		 data0x => SYNTHESIZED_WIRE_28,
		 data1x => SYNTHESIZED_WIRE_29,
		 result => SYNTHESIZED_WIRE_31);


b2v_inst33 : controlunit
PORT MAP(OP => IY_OUT,
		 beq(0) => beq,
		 bgt(0) => bgt,
		 bne(0) => bne,
		 Exop(0) => exop,
		 jump(0) => LOAD_PC,
		 Lmux(0) => LMUX,
		 PC_1(0) => INCR_PC,
		 R_tybe(0) => R_TY,
		 S => SYNTHESIZED_WIRE_46,
		 Smux(0) => HALT,
		 WE(0) => WE);


b2v_inst34 : bit_mux
PORT MAP(sel => R_TY,
		 data0x => IY_OUT(7 DOWNTO 6),
		 data1x => IY_OUT(9 DOWNTO 8),
		 result => SYNTHESIZED_WIRE_4);


SYNTHESIZED_WIRE_37 <= beq AND ZF;


SYNTHESIZED_WIRE_35 <= bgt AND CO;


b2v_inst37 : pc
PORT MAP(clk => SYNTHESIZED_WIRE_54,
		 Reset => reset,
		 LOAD_PC => LOAD_PC,
		 INCR_PC => INCR_PC,
		 Addr_Val_in => SYNTHESIZED_WIRE_31,
		 PC_out => PC_OUT);


SYNTHESIZED_WIRE_29 <= SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_33;


SYNTHESIZED_WIRE_36 <= SYNTHESIZED_WIRE_34 AND bne;


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_35 OR SYNTHESIZED_WIRE_36 OR SYNTHESIZED_WIRE_37;


b2v_inst40 : offset
PORT MAP(in_c => IY_OUT(7 DOWNTO 0),
		 out_c => SYNTHESIZED_WIRE_40);


b2v_inst41 : address
PORT MAP(in_c => IY_OUT,
		 out_c => SYNTHESIZED_WIRE_32);


SYNTHESIZED_WIRE_34 <= NOT(ZF);



b2v_inst43 : lpm_constant1
PORT MAP(		 result => SYNTHESIZED_WIRE_39);


b2v_inst45 : immediate
PORT MAP(in_c => IY_OUT(7 DOWNTO 0),
		 went(0) => exop,
		 out_c => SYNTHESIZED_WIRE_9);


SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_53 AND SYNTHESIZED_WIRE_39;


b2v_inst49 : adder_16bit
PORT MAP(A => SYNTHESIZED_WIRE_40,
		 B => SYNTHESIZED_WIRE_53,
		 Sum => SYNTHESIZED_WIRE_27);


b2v_inst5 : rom0
PORT MAP(clock => SYNTHESIZED_WIRE_42,
		 address => PC_OUT,
		 q => IY_OUT);



b2v_inst51 : adder_16bit
PORT MAP(A => PC_OUT,
		 B => SYNTHESIZED_WIRE_43,
		 Sum => SYNTHESIZED_WIRE_53);


SYNTHESIZED_WIRE_54 <= HALT OR clock;


SYNTHESIZED_WIRE_42 <= NOT(SYNTHESIZED_WIRE_54);



b2v_inst8 : lpm_mux0
PORT MAP(sel => R_TY,
		 data0x => SYNTHESIZED_WIRE_45,
		 data1x => SYNTHESIZED_WIRE_46,
		 result => SYNTHESIZED_WIRE_2);


END bdf_type;